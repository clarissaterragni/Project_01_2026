library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity tb_timer is
    generic (
      clk_freq_hz_g : natural := 100_000_000;
      delay_g       : time    := 2 ms;
      runner_cfg    : string  := ""
    );
end entity tb_timer;

architecture sim of tb_timer is

      constant CLK_PERIOD : time := 1 sec / clk_freq_hz_g;

      signal clk_i   : std_ulogic := '0';
      signal arst_i  : std_ulogic := '0';
      signal start_i : std_ulogic := '0';
      signal done_o  : std_ulogic;

begin
  
      dut : entity work.timer
        generic map (
          clk_freq_hz_g => clk_freq_hz_g,
          delay_g       => delay_g
        )
        port map (
          clk_i   => clk_i,
          arst_i  => arst_i,
          start_i => start_i,
          done_o  => done_o
        );

 
      clk_signal : process begin
          clk_i <= '0';
          wait for CLK_PERIOD / 2;
          clk_i <= '1';
          wait for CLK_PERIOD / 2;
      end process;

  ------------------------------------------------------------------------------
  -- Main test process (VUnit)
  ------------------------------------------------------------------------------
  main : process
      variable t_start : time;
  begin

    test_runner_setup(runner, runner_cfg);

    arst_i <= '1';
    wait for 2 * CLK_PERIOD;
    arst_i <= '0';
    wait for CLK_PERIOD;

    check_equal(done_o, '1', "Timer should be idle after reset");
    
    wait until rising_edge(clk_i);
    start_i <= '1';
    wait until rising_edge(clk_i);
    start_i <= '0';
    wait until rising_edge(clk_i);   -- Had error: added for correct done_o
    
    t_start := now;
    check_equal(done_o, '0', "Timer should be busy after start");

    wait until done_o = '1';


    log("Requested delay: " & time'image(delay_g) & ", Clock frequency: " & integer'image(clk_freq_hz_g) & " Hz" &
        ", Clock period: " & time'image(CLK_PERIOD));

    log("Measured delay (now - t_start): " & time'image(now - t_start));

    if abs((now - t_start) - delay_g) = 0 us then
        log("done_o asserted at EXACT delay");
    else
        log("done_o asserted within one clock period (quantization)");
        check(abs((now - t_start) - delay_g) <= CLK_PERIOD,"done_o asserted within one clock period (quantization)");
    end if;

    -- if correct: get green script when run .py file
    
    log("Test completed successfully");
    
    test_runner_cleanup(runner);

  end process;
end architecture sim;
